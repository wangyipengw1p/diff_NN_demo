/*======================================================
Descripton:


Create:  
Yipeng   wangyipengv@outlook.com  20191127

Modify:

Notes:
1. 

TODO:
=========================================================*/
`include "diff_core_pkg.sv"
